library ieee;
use ieee.std_logic_1164.all;

entity rob is 
    generic(
        size : integer := 256 -- size of the ROB
    );
    port(
        -- INPUTS -------------------------------------------------------------------------------------------
        clk: in std_logic; -- input clock
        clr: in std_logic; -- clear bit
        wr_inst1, wr_inst2: in std_logic; -- write bits for newly decoded instructions 
        wr_ALU1, wr_ALU2: in std_logic; -- write bits for newly executed instructions
        rd: in std_logic; -- read bit for finished instructions
		
        pc_inst1, pc_inst2: in std_logic_vector(15 downto 0); -- PC values for writing the newly decoded instructions
        pc_ALU1, pc_ALU2: in std_logic_vector(15 downto 0); -- PC values for identifying the newly executed instructions
        value_ALU1, value_ALU2: in std_logic_vector(15 downto 0); -- final output values obtained from the execution pipelines
        dest_inst1, dest_inst2: in std_logic_vector(2 downto 0); -- destination registers for newly decoded instructions
        rr1_inst1, rr1_inst2: in std_logic_vector(7 downto 0); -- RR1 for newly decoded instructions
        c_ALU1, z_ALU1, c_ALU2, z_ALU2: in std_logic; -- c and z values obtained from the execution pipelines
        rr2_inst1, rr2_inst2: in std_logic_vector(7 downto 0); -- RR2 for newly decoded instructions
        rr3_inst1, rr3_inst2: in std_logic_vector(7 downto 0); -- RR3 for newly decoded instructions

        -- OUTPUTS -------------------------------------------------------------------------------------------
        rr1_ALU1, rr1_ALU2: out std_logic_vector(7 downto 0); -- RR1 values for both ALU pipelines to which value is written to
        rr2_ALU1, rr2_ALU2, rr3_ALU1, rr3_ALU2: out std_logic_vector(7 downto 0); -- RR2, RR3 values for both ALU pipelines to which flags are written to
        dest_out: out std_logic_vector(2 downto 0); -- destination register for final output
        completed: out std_logic -- bit for when an instruction is completed
	);
end rob;

architecture behavioural of rob is
    -- defining the types required for different-sized columns
    type rob_type_3 is array(size - 1 downto 0) of std_logic_vector(2 downto 0);
    type rob_type_8 is array(size - 1 downto 0) of std_logic_vector(7 downto 0);
    type rob_type_16 is array(size - 1 downto 0) of std_logic_vector(15 downto 0);

    -- defining the required columns, each with (size) entries
    signal rob_pc: rob_type_16:= (others => (others => '0'));
    signal rob_value: rob_type_16:= (others => (others => '0'));

    signal rob_dest: rob_type_3:= (others => (others => '0'));
    signal rob_rr1: rob_type_8:= (others => (others => '0'));

    signal rob_c: std_logic_vector(size - 1 downto 0) := (others => '0');
    signal rob_rr2: rob_type_8:= (others => (others => '0'));

    signal rob_z: std_logic_vector(size - 1 downto 0) := (others => '0');
    signal rob_rr3: rob_type_8:= (others => (others => '0'));

    signal rob_finished: std_logic_vector(size - 1 downto 0) := (others => '0');
    signal rob_completed: std_logic_vector(size - 1 downto 0) := (others => '0');

    -- defining the indexes for read/write, count and the full/empty bits
    signal rd_index, wr_index: integer range 0 to size - 1 := 0;
    signal empty: std_logic := '1';
    signal full: std_logic := '0';
    signal length: integer := 0;

begin
    rob_operation: process(clr, clk) 
        variable count: integer;
        variable head, tail: integer;
        
    begin
        if (clr = '1') then
            -- clear data and indices when reset is set
            rob_pc <= (others => (others => '0'));
            rob_value <= (others => (others => '0'));
            rob_dest <= (others => (others => '0'));
            rob_rr1 <= (others => (others => '0'));
            rob_c <= (others => '0');
            rob_rr2 <= (others => (others => '0'));
            rob_z <= (others => '0');
            rob_rr3 <= (others => (others => '0'));
            rob_finished <= (others => '0');
            rob_completed <= (others => '0');
            wr_index <= 0;
            rd_index <= 0;
            empty <= '1';
            full <= '0';

            count := 0;
            head := 0;
            tail := 0;

        else
            -- FIFO logic and adding newly decoded instructions to the ROB
            if (rising_edge(clk)) then
                -- Writes 1st instruction to the empty entry pointed to by wr_index
                if (wr_inst1 = '1') then
                    rob_pc(tail) <= pc_inst1;
                    rob_dest(tail) <= dest_inst1;
                    rob_rr1(tail) <= rr1_inst1;
                    rob_rr2(tail) <= rr2_inst1;
                    rob_rr3(tail) <= rr3_inst1;
                    rob_finished(tail) <= '0';
                    rob_completed(tail) <= '0';

                    count := count + 1;
                end if;

                -- Write index for the 1st instruction
                if (wr_inst1 = '1' and not (count = size)) then
                    if tail = size - 1 then
                        tail := 0;
                    else
                        tail := tail + 1;
                    end if;
                end if;

                -- Writes 2nd instruction to the empty entry pointed to by wr_index
                if (wr_inst2 = '1') then
                    rob_pc(tail) <= pc_inst2;
                    rob_dest(tail) <= dest_inst2;
                    rob_rr1(tail) <= rr1_inst2;
                    rob_rr2(tail) <= rr2_inst2;
                    rob_rr3(tail) <= rr3_inst2;
                    rob_finished(tail) <= '0';
                    rob_completed(tail) <= '0';

                    count := count + 1;
                end if;

                -- Write index for the 2nd instruction
                if (wr_inst2 = '1' and not (count = size)) then
                    if tail = size - 1 then
                        tail := 0;
                    else
                        tail := tail + 1;
                    end if;
                end if;

                -- Keep track of the rd_index     
                if (rob_finished(i) = '1') then
                    if (rd = '1' and not (count = 0)) then
                        if head = size - 1 then
                            head := 0;
                        else
                            head := head + 1;
                        end if;
    
                        rob_completed(head) <= '1';
                        count := count - 1;
                    end if;
                end if;
                
                -- Writing output values from the execution pipelines
                -- Write executed data from ALU1 into corresponding ROB entry
                if (wr_ALU1 = '1') then
                    for i in 0 to size - 1 loop
                        if (rob_pc(i) = pc_ALU1) then
                            rob_value(i) <= value_ALU1;
                            rob_c(i) <= c_ALU1;
                            rob_z(i) <= z_ALU1;
                            rob_finished(i) <= '1';

                            -- Read rename registers for ALU2 from corresponding ROB entry
                            rr1_ALU1 <= rob_rr1(i);
                            rr2_ALU1 <= rob_rr2(i);
                            rr3_ALU1 <= rob_rr3(i);
                            exit;
                        end if;
                    end loop;

                else
                    rr1_ALU1 <= (others => '0');
                    rr2_ALU1 <= (others => '0');
                    rr3_ALU1 <= (others => '0');
                end if;

                -- Write executed data from ALU2 into corresponding ROB entry
                if (wr_ALU2 = '1') then
                    for i in 0 to size-1 loop
                        if (rob_pc(i) = pc_ALU2) then
                            rob_value(i) <= value_ALU2;
                            rob_c(i) <= c_ALU2;
                            rob_z(i) <= z_ALU2;
                            rob_finished(i) <= '1';

                            -- Read rename registers for ALU2 from corresponding ROB entry
                            rr1_ALU2 <= rob_rr1(i);
                            rr2_ALU2 <= rob_rr2(i);
                            rr3_ALU2 <= rob_rr3(i);
                            exit;
                        end if;
                    end loop;

                else
                    rr1_ALU2 <= (others => '0');
                    rr2_ALU2 <= (others => '0');
                    rr3_ALU2 <= (others => '0');
                end if;
            end if;

            rd_index <= head;
            wr_index <= tail;
            length <= count;

            -- Check empty, full
            if (count = 0) then
                empty <= '1';
            else
                empty <= '0';
            end if;

            if (count = size) then
                full <= '1';
            else
                full <= '0';
            end if;
        end if;
    end process rob_operation;

    -- Value from entry pointed to by rd_index
    dest_out <= rob_dest(rd_index);
    completed <= rob_completed(rd_index);
end architecture behavioural;